module inverter(out, in);
  output out;
  input in;
  assign out = ~in;
endmodule
