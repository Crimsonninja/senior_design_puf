module puf_1_bit(en32, );
  output [8:0]
  input [32:0] en32;

  shift_register SR();

endmodule
